`timescale 1ns / 1ps

/// @brief 5到32位译码器
module Decoder5T32(
    input [4: 0] DataIn,
    input Enable,
    output reg [31: 0]Y);

    always@(Enable or DataIn) begin
        if(Enable) begin
            case(DataIn)
                5'b00000 : Y <= 32'b00000000000000000000000000000001;
                5'b00001 : Y <= 32'b00000000000000000000000000000010;
                5'b00010 : Y <= 32'b00000000000000000000000000000100;
                5'b00011 : Y <= 32'b00000000000000000000000000001000;
                5'b00100 : Y <= 32'b00000000000000000000000000010000;
                5'b00101 : Y <= 32'b00000000000000000000000000100000;
                5'b00110 : Y <= 32'b00000000000000000000000001000000;
                5'b00111 : Y <= 32'b00000000000000000000000010000000;
                5'b01000 : Y <= 32'b00000000000000000000000100000000;
                5'b01001 : Y <= 32'b00000000000000000000001000000000;
                5'b01010 : Y <= 32'b00000000000000000000010000000000;
                5'b01011 : Y <= 32'b00000000000000000000100000000000;
                5'b01100 : Y <= 32'b00000000000000000001000000000000;
                5'b01101 : Y <= 32'b00000000000000000010000000000000;
                5'b01110 : Y <= 32'b00000000000000000100000000000000;
                5'b01111 : Y <= 32'b00000000000000001000000000000000;
                5'b10000 : Y <= 32'b00000000000000010000000000000000;
                5'b10001 : Y <= 32'b00000000000000100000000000000000;
                5'b10010 : Y <= 32'b00000000000001000000000000000000;
                5'b10011 : Y <= 32'b00000000000010000000000000000000;
                5'b10100 : Y <= 32'b00000000000100000000000000000000;
                5'b10101 : Y <= 32'b00000000001000000000000000000000;
                5'b10110 : Y <= 32'b00000000010000000000000000000000;
                5'b10111 : Y <= 32'b00000000100000000000000000000000;
                5'b11000 : Y <= 32'b00000001000000000000000000000000;
                5'b11001 : Y <= 32'b00000010000000000000000000000000;
                5'b11010 : Y <= 32'b00000100000000000000000000000000;
                5'b11011 : Y <= 32'b00001000000000000000000000000000;
                5'b11100 : Y <= 32'b00010000000000000000000000000000;
                5'b11101 : Y <= 32'b00100000000000000000000000000000;
                5'b11110 : Y <= 32'b01000000000000000000000000000000;
                5'b11111 : Y <= 32'b10000000000000000000000000000000;
            endcase
        end 
        else Y <= 32'b00000000000000000000000000000000;
    end
endmodule
